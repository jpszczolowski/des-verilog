module S8(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 13 :
          (in == 1) ? 1 :
          (in == 2) ? 2 :
          (in == 3) ? 15 :
          (in == 4) ? 8 :
          (in == 5) ? 13 :
          (in == 6) ? 4 :
          (in == 7) ? 8 :
          (in == 8) ? 6 :
          (in == 9) ? 10 :
          (in == 10) ? 15 :
          (in == 11) ? 3 :
          (in == 12) ? 11 :
          (in == 13) ? 7 :
          (in == 14) ? 1 :
          (in == 15) ? 4 :
          (in == 16) ? 10 :
          (in == 17) ? 12 :
          (in == 18) ? 9 :
          (in == 19) ? 5 :
          (in == 20) ? 3 :
          (in == 21) ? 6 :
          (in == 22) ? 14 :
          (in == 23) ? 11 :
          (in == 24) ? 5 :
          (in == 25) ? 0 :
          (in == 26) ? 0 :
          (in == 27) ? 14 :
          (in == 28) ? 12 :
          (in == 29) ? 9 :
          (in == 30) ? 7 :
          (in == 31) ? 2 :
          (in == 32) ? 7 :
          (in == 33) ? 2 :
          (in == 34) ? 11 :
          (in == 35) ? 1 :
          (in == 36) ? 4 :
          (in == 37) ? 14 :
          (in == 38) ? 1 :
          (in == 39) ? 7 :
          (in == 40) ? 9 :
          (in == 41) ? 4 :
          (in == 42) ? 12 :
          (in == 43) ? 10 :
          (in == 44) ? 14 :
          (in == 45) ? 8 :
          (in == 46) ? 2 :
          (in == 47) ? 13 :
          (in == 48) ? 0 :
          (in == 49) ? 15 :
          (in == 50) ? 6 :
          (in == 51) ? 12 :
          (in == 52) ? 10 :
          (in == 53) ? 9 :
          (in == 54) ? 13 :
          (in == 55) ? 0 :
          (in == 56) ? 15 :
          (in == 57) ? 3 :
          (in == 58) ? 3 :
          (in == 59) ? 5 :
          (in == 60) ? 5 :
          (in == 61) ? 6 :
          (in == 62) ? 8 :
          (in == 63) ? 11 :
          0;
endmodule
