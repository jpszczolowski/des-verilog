module S1(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 14 :
          (in == 1) ? 0 :
          (in == 2) ? 4 :
          (in == 3) ? 15 :
          (in == 4) ? 13 :
          (in == 5) ? 7 :
          (in == 6) ? 1 :
          (in == 7) ? 4 :
          (in == 8) ? 2 :
          (in == 9) ? 14 :
          (in == 10) ? 15 :
          (in == 11) ? 2 :
          (in == 12) ? 11 :
          (in == 13) ? 13 :
          (in == 14) ? 8 :
          (in == 15) ? 1 :
          (in == 16) ? 3 :
          (in == 17) ? 10 :
          (in == 18) ? 10 :
          (in == 19) ? 6 :
          (in == 20) ? 6 :
          (in == 21) ? 12 :
          (in == 22) ? 12 :
          (in == 23) ? 11 :
          (in == 24) ? 5 :
          (in == 25) ? 9 :
          (in == 26) ? 9 :
          (in == 27) ? 5 :
          (in == 28) ? 0 :
          (in == 29) ? 3 :
          (in == 30) ? 7 :
          (in == 31) ? 8 :
          (in == 32) ? 4 :
          (in == 33) ? 15 :
          (in == 34) ? 1 :
          (in == 35) ? 12 :
          (in == 36) ? 14 :
          (in == 37) ? 8 :
          (in == 38) ? 8 :
          (in == 39) ? 2 :
          (in == 40) ? 13 :
          (in == 41) ? 4 :
          (in == 42) ? 6 :
          (in == 43) ? 9 :
          (in == 44) ? 2 :
          (in == 45) ? 1 :
          (in == 46) ? 11 :
          (in == 47) ? 7 :
          (in == 48) ? 15 :
          (in == 49) ? 5 :
          (in == 50) ? 12 :
          (in == 51) ? 11 :
          (in == 52) ? 9 :
          (in == 53) ? 3 :
          (in == 54) ? 7 :
          (in == 55) ? 14 :
          (in == 56) ? 3 :
          (in == 57) ? 10 :
          (in == 58) ? 10 :
          (in == 59) ? 0 :
          (in == 60) ? 5 :
          (in == 61) ? 6 :
          (in == 62) ? 0 :
          (in == 63) ? 13 :
          0;
endmodule
