module S6(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 12 :
          (in == 1) ? 10 :
          (in == 2) ? 1 :
          (in == 3) ? 15 :
          (in == 4) ? 10 :
          (in == 5) ? 4 :
          (in == 6) ? 15 :
          (in == 7) ? 2 :
          (in == 8) ? 9 :
          (in == 9) ? 7 :
          (in == 10) ? 2 :
          (in == 11) ? 12 :
          (in == 12) ? 6 :
          (in == 13) ? 9 :
          (in == 14) ? 8 :
          (in == 15) ? 5 :
          (in == 16) ? 0 :
          (in == 17) ? 6 :
          (in == 18) ? 13 :
          (in == 19) ? 1 :
          (in == 20) ? 3 :
          (in == 21) ? 13 :
          (in == 22) ? 4 :
          (in == 23) ? 14 :
          (in == 24) ? 14 :
          (in == 25) ? 0 :
          (in == 26) ? 7 :
          (in == 27) ? 11 :
          (in == 28) ? 5 :
          (in == 29) ? 3 :
          (in == 30) ? 11 :
          (in == 31) ? 8 :
          (in == 32) ? 9 :
          (in == 33) ? 4 :
          (in == 34) ? 14 :
          (in == 35) ? 3 :
          (in == 36) ? 15 :
          (in == 37) ? 2 :
          (in == 38) ? 5 :
          (in == 39) ? 12 :
          (in == 40) ? 2 :
          (in == 41) ? 9 :
          (in == 42) ? 8 :
          (in == 43) ? 5 :
          (in == 44) ? 12 :
          (in == 45) ? 15 :
          (in == 46) ? 3 :
          (in == 47) ? 10 :
          (in == 48) ? 7 :
          (in == 49) ? 11 :
          (in == 50) ? 0 :
          (in == 51) ? 14 :
          (in == 52) ? 4 :
          (in == 53) ? 1 :
          (in == 54) ? 10 :
          (in == 55) ? 7 :
          (in == 56) ? 1 :
          (in == 57) ? 6 :
          (in == 58) ? 13 :
          (in == 59) ? 0 :
          (in == 60) ? 11 :
          (in == 61) ? 8 :
          (in == 62) ? 6 :
          (in == 63) ? 13 :
          0;
endmodule
