module S4(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 7 :
          (in == 1) ? 13 :
          (in == 2) ? 13 :
          (in == 3) ? 8 :
          (in == 4) ? 14 :
          (in == 5) ? 11 :
          (in == 6) ? 3 :
          (in == 7) ? 5 :
          (in == 8) ? 0 :
          (in == 9) ? 6 :
          (in == 10) ? 6 :
          (in == 11) ? 15 :
          (in == 12) ? 9 :
          (in == 13) ? 0 :
          (in == 14) ? 10 :
          (in == 15) ? 3 :
          (in == 16) ? 1 :
          (in == 17) ? 4 :
          (in == 18) ? 2 :
          (in == 19) ? 7 :
          (in == 20) ? 8 :
          (in == 21) ? 2 :
          (in == 22) ? 5 :
          (in == 23) ? 12 :
          (in == 24) ? 11 :
          (in == 25) ? 1 :
          (in == 26) ? 12 :
          (in == 27) ? 10 :
          (in == 28) ? 4 :
          (in == 29) ? 14 :
          (in == 30) ? 15 :
          (in == 31) ? 9 :
          (in == 32) ? 10 :
          (in == 33) ? 3 :
          (in == 34) ? 6 :
          (in == 35) ? 15 :
          (in == 36) ? 9 :
          (in == 37) ? 0 :
          (in == 38) ? 0 :
          (in == 39) ? 6 :
          (in == 40) ? 12 :
          (in == 41) ? 10 :
          (in == 42) ? 11 :
          (in == 43) ? 1 :
          (in == 44) ? 7 :
          (in == 45) ? 13 :
          (in == 46) ? 13 :
          (in == 47) ? 8 :
          (in == 48) ? 15 :
          (in == 49) ? 9 :
          (in == 50) ? 1 :
          (in == 51) ? 4 :
          (in == 52) ? 3 :
          (in == 53) ? 5 :
          (in == 54) ? 14 :
          (in == 55) ? 11 :
          (in == 56) ? 5 :
          (in == 57) ? 12 :
          (in == 58) ? 2 :
          (in == 59) ? 7 :
          (in == 60) ? 8 :
          (in == 61) ? 2 :
          (in == 62) ? 4 :
          (in == 63) ? 14 :
          0;
endmodule
