module S3(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 10 :
          (in == 1) ? 13 :
          (in == 2) ? 0 :
          (in == 3) ? 7 :
          (in == 4) ? 9 :
          (in == 5) ? 0 :
          (in == 6) ? 14 :
          (in == 7) ? 9 :
          (in == 8) ? 6 :
          (in == 9) ? 3 :
          (in == 10) ? 3 :
          (in == 11) ? 4 :
          (in == 12) ? 15 :
          (in == 13) ? 6 :
          (in == 14) ? 5 :
          (in == 15) ? 10 :
          (in == 16) ? 1 :
          (in == 17) ? 2 :
          (in == 18) ? 13 :
          (in == 19) ? 8 :
          (in == 20) ? 12 :
          (in == 21) ? 5 :
          (in == 22) ? 7 :
          (in == 23) ? 14 :
          (in == 24) ? 11 :
          (in == 25) ? 12 :
          (in == 26) ? 4 :
          (in == 27) ? 11 :
          (in == 28) ? 2 :
          (in == 29) ? 15 :
          (in == 30) ? 8 :
          (in == 31) ? 1 :
          (in == 32) ? 13 :
          (in == 33) ? 1 :
          (in == 34) ? 6 :
          (in == 35) ? 10 :
          (in == 36) ? 4 :
          (in == 37) ? 13 :
          (in == 38) ? 9 :
          (in == 39) ? 0 :
          (in == 40) ? 8 :
          (in == 41) ? 6 :
          (in == 42) ? 15 :
          (in == 43) ? 9 :
          (in == 44) ? 3 :
          (in == 45) ? 8 :
          (in == 46) ? 0 :
          (in == 47) ? 7 :
          (in == 48) ? 11 :
          (in == 49) ? 4 :
          (in == 50) ? 1 :
          (in == 51) ? 15 :
          (in == 52) ? 2 :
          (in == 53) ? 14 :
          (in == 54) ? 12 :
          (in == 55) ? 3 :
          (in == 56) ? 5 :
          (in == 57) ? 11 :
          (in == 58) ? 10 :
          (in == 59) ? 5 :
          (in == 60) ? 14 :
          (in == 61) ? 2 :
          (in == 62) ? 7 :
          (in == 63) ? 12 :
          0;
endmodule
