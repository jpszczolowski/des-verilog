module S2(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 15 :
          (in == 1) ? 3 :
          (in == 2) ? 1 :
          (in == 3) ? 13 :
          (in == 4) ? 8 :
          (in == 5) ? 4 :
          (in == 6) ? 14 :
          (in == 7) ? 7 :
          (in == 8) ? 6 :
          (in == 9) ? 15 :
          (in == 10) ? 11 :
          (in == 11) ? 2 :
          (in == 12) ? 3 :
          (in == 13) ? 8 :
          (in == 14) ? 4 :
          (in == 15) ? 14 :
          (in == 16) ? 9 :
          (in == 17) ? 12 :
          (in == 18) ? 7 :
          (in == 19) ? 0 :
          (in == 20) ? 2 :
          (in == 21) ? 1 :
          (in == 22) ? 13 :
          (in == 23) ? 10 :
          (in == 24) ? 12 :
          (in == 25) ? 6 :
          (in == 26) ? 0 :
          (in == 27) ? 9 :
          (in == 28) ? 5 :
          (in == 29) ? 11 :
          (in == 30) ? 10 :
          (in == 31) ? 5 :
          (in == 32) ? 0 :
          (in == 33) ? 13 :
          (in == 34) ? 14 :
          (in == 35) ? 8 :
          (in == 36) ? 7 :
          (in == 37) ? 10 :
          (in == 38) ? 11 :
          (in == 39) ? 1 :
          (in == 40) ? 10 :
          (in == 41) ? 3 :
          (in == 42) ? 4 :
          (in == 43) ? 15 :
          (in == 44) ? 13 :
          (in == 45) ? 4 :
          (in == 46) ? 1 :
          (in == 47) ? 2 :
          (in == 48) ? 5 :
          (in == 49) ? 11 :
          (in == 50) ? 8 :
          (in == 51) ? 6 :
          (in == 52) ? 12 :
          (in == 53) ? 7 :
          (in == 54) ? 6 :
          (in == 55) ? 12 :
          (in == 56) ? 9 :
          (in == 57) ? 0 :
          (in == 58) ? 3 :
          (in == 59) ? 5 :
          (in == 60) ? 2 :
          (in == 61) ? 14 :
          (in == 62) ? 15 :
          (in == 63) ? 9 :
          0;
endmodule
