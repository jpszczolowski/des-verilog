module S7(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 4 :
          (in == 1) ? 13 :
          (in == 2) ? 11 :
          (in == 3) ? 0 :
          (in == 4) ? 2 :
          (in == 5) ? 11 :
          (in == 6) ? 14 :
          (in == 7) ? 7 :
          (in == 8) ? 15 :
          (in == 9) ? 4 :
          (in == 10) ? 0 :
          (in == 11) ? 9 :
          (in == 12) ? 8 :
          (in == 13) ? 1 :
          (in == 14) ? 13 :
          (in == 15) ? 10 :
          (in == 16) ? 3 :
          (in == 17) ? 14 :
          (in == 18) ? 12 :
          (in == 19) ? 3 :
          (in == 20) ? 9 :
          (in == 21) ? 5 :
          (in == 22) ? 7 :
          (in == 23) ? 12 :
          (in == 24) ? 5 :
          (in == 25) ? 2 :
          (in == 26) ? 10 :
          (in == 27) ? 15 :
          (in == 28) ? 6 :
          (in == 29) ? 8 :
          (in == 30) ? 1 :
          (in == 31) ? 6 :
          (in == 32) ? 1 :
          (in == 33) ? 6 :
          (in == 34) ? 4 :
          (in == 35) ? 11 :
          (in == 36) ? 11 :
          (in == 37) ? 13 :
          (in == 38) ? 13 :
          (in == 39) ? 8 :
          (in == 40) ? 12 :
          (in == 41) ? 1 :
          (in == 42) ? 3 :
          (in == 43) ? 4 :
          (in == 44) ? 7 :
          (in == 45) ? 10 :
          (in == 46) ? 14 :
          (in == 47) ? 7 :
          (in == 48) ? 10 :
          (in == 49) ? 9 :
          (in == 50) ? 15 :
          (in == 51) ? 5 :
          (in == 52) ? 6 :
          (in == 53) ? 0 :
          (in == 54) ? 8 :
          (in == 55) ? 15 :
          (in == 56) ? 0 :
          (in == 57) ? 14 :
          (in == 58) ? 5 :
          (in == 59) ? 2 :
          (in == 60) ? 9 :
          (in == 61) ? 3 :
          (in == 62) ? 2 :
          (in == 63) ? 12 :
          0;
endmodule
