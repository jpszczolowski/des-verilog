module S5(input [6:1] in, output [4:1] out);
  assign out =
          (in == 0) ? 2 :
          (in == 1) ? 14 :
          (in == 2) ? 12 :
          (in == 3) ? 11 :
          (in == 4) ? 4 :
          (in == 5) ? 2 :
          (in == 6) ? 1 :
          (in == 7) ? 12 :
          (in == 8) ? 7 :
          (in == 9) ? 4 :
          (in == 10) ? 10 :
          (in == 11) ? 7 :
          (in == 12) ? 11 :
          (in == 13) ? 13 :
          (in == 14) ? 6 :
          (in == 15) ? 1 :
          (in == 16) ? 8 :
          (in == 17) ? 5 :
          (in == 18) ? 5 :
          (in == 19) ? 0 :
          (in == 20) ? 3 :
          (in == 21) ? 15 :
          (in == 22) ? 15 :
          (in == 23) ? 10 :
          (in == 24) ? 13 :
          (in == 25) ? 3 :
          (in == 26) ? 0 :
          (in == 27) ? 9 :
          (in == 28) ? 14 :
          (in == 29) ? 8 :
          (in == 30) ? 9 :
          (in == 31) ? 6 :
          (in == 32) ? 4 :
          (in == 33) ? 11 :
          (in == 34) ? 2 :
          (in == 35) ? 8 :
          (in == 36) ? 1 :
          (in == 37) ? 12 :
          (in == 38) ? 11 :
          (in == 39) ? 7 :
          (in == 40) ? 10 :
          (in == 41) ? 1 :
          (in == 42) ? 13 :
          (in == 43) ? 14 :
          (in == 44) ? 7 :
          (in == 45) ? 2 :
          (in == 46) ? 8 :
          (in == 47) ? 13 :
          (in == 48) ? 15 :
          (in == 49) ? 6 :
          (in == 50) ? 9 :
          (in == 51) ? 15 :
          (in == 52) ? 12 :
          (in == 53) ? 0 :
          (in == 54) ? 5 :
          (in == 55) ? 9 :
          (in == 56) ? 6 :
          (in == 57) ? 10 :
          (in == 58) ? 3 :
          (in == 59) ? 4 :
          (in == 60) ? 0 :
          (in == 61) ? 5 :
          (in == 62) ? 14 :
          (in == 63) ? 3 :
          0;
endmodule
